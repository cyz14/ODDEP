library IEEE;USE IEEE.STD_LOGIC_1164.ALL;USE IEEE.STD_LOGIC_ARITH.ALL;USE IEEE.STD_LOGIC_UNSIGNED.ALL;entity digitalEO is    port(        oe:in STD_LOGIC;        six6:out STD_LOGIC;        six7:out STD_LOGIC;        egt8:out STD_LOGIC;        egt9:out STD_LOGIC;        eiA:out STD_LOGIC;        eiB:out STD_LOGIC        );end entity;architecture eo_digital of digitalEO isbegin    six6 <= not oe;    egt8 <= not oe;    eiA <= not oe;    six7 <= oe;    egt9 <= oe;    eiB <= oe;end eo_digital;